`ifndef MEMORY_ACCESS_VH_
`define MEMORY_ACCESS_VH_

`define ACC_WORD 2'b00
`define ACC_DWORD 2'b01
`define ACC_BURST 2'b10

`endif // MEMORY_ACCESS_VH_
