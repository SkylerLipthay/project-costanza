`ifndef REGISTERS_VH_
`define REGISTERS_VH_

`define REG_A 4'd0
`define REG_B 4'd1
`define REG_C 4'd2
`define REG_D 4'd3
`define REG_E 4'd4
`define REG_F 4'd5
`define REG_MH 4'd6
`define REG_ML 4'd7
`define REG_J1 4'd8
`define REG_J2 4'd9
`define REG_G 4'd10
`define REG_H 4'd11
`define REG_X 4'd12
`define REG_Y 4'd13
`define REG_0 4'd14
`define REG_1 4'd15

`endif // REGISTERS_VH_
