`ifndef INSTRUCTIONS_VH_
`define INSTRUCTIONS_VH_

`define INS_MOV_REG 8'b00000000
`define INS_MOV_LIT 8'b00000001
`define INS_LD 8'b00000010
`define INS_ST 8'b00000011
`define INS_LEA 8'b00000100
`define INS_BR 8'b00010000
`define INS_BRL 8'b00010001
`define INS_BRLE 8'b00010010
`define INS_BRG 8'b00010011
`define INS_BRGE 8'b00010100
`define INS_BRE 8'b00010101
`define INS_BRNE 8'b00010110
`define INS_BRB 8'b00010111
`define INS_BRBE 8'b00011000
`define INS_BRA 8'b00011001
`define INS_BRAE 8'b00011010
`define INS_ADD 8'b00110000
`define INS_SUB 8'b00110001
`define INS_AND 8'b00110010
`define INS_OR 8'b00110011
`define INS_XOR 8'b00110100
`define INS_NOT 8'b00110101
`define INS_CMP 8'b00110110
`define INS_SHL 8'b00110111
`define INS_SHR 8'b00111000
`define INS_RL 8'b00111001
`define INS_RR 8'b00111010
`define INS_NEG 8'b00111011
`define INS_ADDMA 8'b01110100
`define INS_SUBMA 8'b01110101
`define INS_SSP 8'b01000000
`define INS_PUSH 8'b01000001
`define INS_POP 8'b01000010
`define INS_CALL 8'b01000101
`define INS_RET 8'b01000110
`define INS_LSP 8'b01000111
`define INS_NOP 8'b01010000
`define INS_HALT 8'b01010001
`define INS_HRD 8'b01010010
`define INS_HWR 8'b01010011
`define INS_SNDA 8'b01010100
`define INS_SNDL 8'b01010101
`define INS_SNDR 8'b01010110
`define INS_SNDW 8'b01010111
`define INS_SNDP 8'b01011000
`define INS_IMGD 8'b01011001
`define INS_IMGCD 8'b01011010
`define INS_IMGC 8'b01011011
`define INS_IMGA 8'b01011100
`define INS_FLIP 8'b01011101

`endif // INSTRUCTIONS_VH_
